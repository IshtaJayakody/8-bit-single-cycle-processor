/*
Module  : Data Cache 
Author  : Isuru Nawinne, Kisaru Liyanage
Date    : 25/05/2020

Description	:

This file presents a skeleton implementation of the cache controller using a Finite State Machine model. Note that this code is not complete.
*/

`timescale 1ns/100ps

module dcache (
    clock,
    reset,
    read,
    write,
    address,
    writedata,
    readdata,
    busywait,
    mem_busywait,
    mem_read,
    mem_write,
    mem_writedata,
    mem_readdata,
    mem_address
);
    //This is the module for cache memory
    //Here is the port declaration
    input clock, reset,read,write; // Initially clock, reset, read, write signals defined as inputs 
    output reg busywait; // Then the busywait signal is defined as reg type because it is a control signal
    input [7:0] writedata, address; // writedata and address are 8-bit inputs
    output reg [7:0] readdata; // readdata is defined as a 8-bit output  
    input mem_busywait; // Then mem_busywait signal is declared as a input which generated by the data memory
    output reg mem_read; // mem_read, mem_write signals are outputs which are controlling the data memory. So the define as output reg type 
    output reg mem_write;
    output reg [31:0] mem_writedata; // mem_writedata and mem_readdata are 32-bit wires
    input [31:0] mem_readdata;
    output reg [5:0] mem_address; // mem_address is a output which carries 5-bit address to the data memeory

    wire valid_bit, dirty, hit; // Then dirty, hit and valid_bit ara defined as wires 
    wire [2:0] tag, index; // tan and index are 3-bit wires
    reg [7:0] word_selector; // This word_selector is use for read data according to the offset of the address

    ///////////////////////////////
    reg [36:0] cacheMem_array [7:0]; // Finally here we are defining 8 memory blocks in the cache memory 
    //extra 5 bits for validbot =1 , dirtybit = 1 , tag=3
    

    /*
    Combinational part for indexing, tag comparison for hit deciding, etc.
    ...
    ...
    */

    // Initially, after arriving a new address to the memory dirty bit, valid_bit, index and tag are extracted after 1 time unit delay
    assign #1 index = address[4:2];
    assign #1 valid_bit =  cacheMem_array[address[4:2]][35];
    assign #1 dirty = cacheMem_array[address[4:2]][36];
    assign #1 tag = cacheMem_array[address[4:2]][34:32];

    // Then hit signal is generated considering valid bit, tag of the existing meory block and tag part of the address.
    //This takes 0.9 time unit delay
    assign #0.9 hit = ((tag == address[7:5])&& valid_bit) ? 1'b1 : 1'b0;

    // This always block is used to output the data which a stored in cache to the register file
    // Always block is sensitive to address, hit, read and write
    always @ (address, hit,read,write)
    begin
        // If there is a read and a hit, initially word selecter is updated in 1 time unit according to the offset
        if(read && hit)
        begin
            case (address[1:0])
                2'b00: #1 word_selector = cacheMem_array[address[4:2]][7:0];
                2'b01: #1 word_selector = cacheMem_array[address[4:2]][15:8];
                2'b10: #1 word_selector = cacheMem_array[address[4:2]][23:16];
                2'b11: #1 word_selector = cacheMem_array[address[4:2]][31:24];
            endcase
            // Then assign that value to readdata
            readdata = word_selector;
        end
    end

    // This always block is used to update the cache when there is a writing operation
    // always block is sensitive to hit
    always @ (hit)
    begin
        //If there is a wtite and a hit, initially cache memory is updated according to the offset. This takes dalay of 1 time unit
        if(write && hit)
        begin
            case (address[1:0])
                2'b00: #1 cacheMem_array[address[4:2]][7:0] = writedata;
                2'b01: #1 cacheMem_array[address[4:2]][15:8] = writedata;
                2'b10: #1 cacheMem_array[address[4:2]][23:16] = writedata;
                2'b11: #1 cacheMem_array[address[4:2]][31:24] = writedata;
            endcase
            //Finally dirty bit is updated
            cacheMem_array[address[4:2]][36] = 1;
        end
    end

    // This always block is used to update cache from the data memory
    // always block is sensitive to mem_read
    always @ ( mem_read)
    begin
        // If mem_read equals to zero followig set of code will be triggered after 1 time unit delay
        if(mem_read == 0)
        begin
            #1
            cacheMem_array[address[4:2]][36] = 0; // Initially dirty bit is set as 0
            cacheMem_array[address[4:2]][35] = 1; // then valid bit is set as 1
            cacheMem_array[address[4:2]][34:32] = address[7:5]; // then the tag part of the cache memory block is set 
            cacheMem_array[address[4:2]][31:0] = mem_readdata;// finally read data from memory will assign to the correspondig cache memory block
        end
    end

    
    /* Cache Controller FSM Start */

    parameter IDLE = 3'b000, MEM_READ = 3'b001, MEM_WRITE = 3'b010;
    reg [2:0] state, next_state;

    // Here is combinational next state logic
    always @(*)
    begin
        case (state)
            IDLE:
                // In the ideal state if there is a read or write operation and dirty bit and hit equals to zero 
                //next state is assigned as MEM_READ
                if ((read || write) && !dirty && !hit)  
                    next_state = MEM_READ;
                //if there is a read or write operation and dirty bit is 1 and there is a miss next state is assigned as MEM_WRITE
                else if ((read || write) && dirty && !hit)
                    next_state = MEM_WRITE;
                // Otherwise it remains in ideal state
                else
                    next_state = IDLE;
            
            MEM_READ:
                // In the memory reading state if mem_busywait signal is 0, next state is assigned as ideal
                if (!mem_busywait)
                    next_state = IDLE;
                // Otherwise it remains in memory reading state 
                else    
                    next_state = MEM_READ;
            MEM_WRITE:
                // In the memory writing state if mem_busywait signal is 0, next state is assigned as MEM_READ
                if (!mem_busywait)
                    next_state = MEM_READ;
                // Otherwise it remains in memory writing state 
                else
                    next_state = MEM_WRITE;
        endcase
    end

    // Here is the combinational output logic
    // This always block is triggered to all the changes in the cache while simulating
    always @(*)
    begin
        case(state)
            IDLE:
            begin
                mem_read = 0;
                mem_write = 0;
                mem_address = 8'dx;
                mem_writedata = 32'dx;
                if((read || write) && !hit) // if there is a read or wtire opearation and there is miss busywait is assigned as 1
                    busywait = 1;
                else
                    busywait = 0;
            end
         
            MEM_READ: 
            begin
                mem_read = 1;
                mem_write = 0;
                mem_address = {address[7:5], index};
                mem_writedata = 32'dx;
                busywait = 1;
            end

            MEM_WRITE:
            begin
                mem_read = 0;
                mem_write = 1;
                mem_address = {cacheMem_array[address[4:2]][34:32], index};
                mem_writedata = cacheMem_array[address[4:2]][31:0];
                busywait = 1;
            end
            
        endcase
    end

    // Here is sequential logic for state transitioning and reset the cache memory
    integer i; 
    always @(posedge clock, reset)
    begin
        // If reset signal is high, state is initialized to the ideal state. And all the cache memory data is cleared
        if(reset)
        begin
            state = IDLE;
            for (i=0;i<8; i=i+1)
            begin
            cacheMem_array[i] = 0;
            end
        end
        else
        // Otherwise circuit will be moved to next state.
        begin
            state = next_state;
        end
    end

    /* Cache Controller FSM End */

endmodule